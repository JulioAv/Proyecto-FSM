module testbench();
reg clock, reset, V0, V1, V2, B0, B1, B2, P0, P1, P2, P3;
wire V0o, V1o, V2o, B0o, B1o, B2o;

FSM f1(clock, reset, V0, V1, V2, B0, B1, B2, P0, P1, P2, P3, V0o, V1o, V2o, B0o, B1o, B2o);
always
	#1 clock <=~clock;
	
	initial begin
	#1
	$display("Control de Volumen y Bajo");
	$display("V2  V1  V0  B2  B1  B0  P3  P2  P1  P0 | V2o  V1o  V0o  B2o  B1o  B0o");
	$display("---------------------------------------|-----------------------------");
	$monitor("%b  %b  %b  %b  %b  %b  %b  %b  %b  %b  |  %b  %b  %b  %b  %b  %b", V2, V1, V0, B2, B1, B0, P3, P2, P1, P0, V2o, V1o, V0o, B2o, B1o, B0);
	end
	initial begin
		reset=0; clock=0;
	#1 V2=0; V1=0; V0=0; B2=0; B1=0; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=0; V0=1; B2=0; B1=0; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=1; V0=0; B2=0; B1=0; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=1; V0=1; B2=0; B1=0; B0=0; P3=0; P2=0; P1=0; P0=0;
	
	#1 V2=0; V1=0; V0=0; B2=0; B1=0; B0=1; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=0; V0=0; B2=0; B1=1; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=0; V0=0; B2=0; B1=1; B0=1; P3=0; P2=0; P1=0; P0=0;
	
	#1 V2=0; V1=0; V0=1; B2=0; B1=0; B0=1; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=0; V0=1; B2=0; B1=1; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=0; V0=1; B2=0; B1=1; B0=1; P3=0; P2=0; P1=0; P0=0;
	
	#1 V2=0; V1=1; V0=0; B2=0; B1=0; B0=1; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=1; V0=0; B2=0; B1=1; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=1; V0=0; B2=0; B1=1; B0=1; P3=0; P2=0; P1=0; P0=0;
	
	#1 V2=0; V1=1; V0=1; B2=0; B1=0; B0=1; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=1; V0=1; B2=0; B1=1; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=1; V0=1; B2=0; B1=1; B0=1; P3=0; P2=0; P1=0; P0=0;
	
	#1 V2=0; V1=0; V0=1; B2=0; B1=0; B0=1; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=0; V0=1; B2=0; B1=1; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=0; V0=1; B2=0; B1=1; B0=1; P3=0; P2=0; P1=0; P0=0;
	
	#1 V2=0; V1=1; V0=1; B2=0; B1=0; B0=1; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=1; V0=1; B2=0; B1=1; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=1; V0=1; B2=0; B1=1; B0=1; P3=0; P2=0; P1=0; P0=0;

	
	#1 V2=1; V1=0; V0=0; B2=0; B1=0; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=1; V1=0; V0=0; B2=0; B1=0; B0=1; P3=0; P2=0; P1=0; P0=0;
	#1 V2=1; V1=0; V0=0; B2=0; B1=1; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=1; V1=0; V0=0; B2=0; B1=1; B0=1; P3=0; P2=0; P1=0; P0=0;	
	
	#1 V2=0; V1=0; V0=0; B2=1; B1=0; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=0; V0=1; B2=1; B1=0; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=1; V0=0; B2=1; B1=0; B0=0; P3=0; P2=0; P1=0; P0=0;
	#1 V2=0; V1=1; V0=1; B2=1; B1=0; B0=0; P3=0; P2=0; P1=0; P0=0;	
	
	#1 V2=0; V1=0; V0=0; B2=0; B1=0; B0=0; P3=0; P2=0; P1=0; P0=1;
	#1 V2=0; V1=0; V0=0; B2=0; B1=0; B0=0; P3=0; P2=0; P1=1; P0=0;
	#1 V2=0; V1=0; V0=0; B2=0; B1=0; B0=0; P3=0; P2=0; P1=1; P0=1;
	#1 V2=0; V1=0; V0=0; B2=0; B1=0; B0=0; P3=0; P2=1; P1=0; P0=0;	
	#1 V2=0; V1=0; V0=0; B2=0; B1=0; B0=0; P3=0; P2=1; P1=0; P0=1;
	#1 V2=0; V1=0; V0=0; B2=0; B1=0; B0=0; P3=0; P2=1; P1=1; P0=0;
	#1 V2=0; V1=0; V0=0; B2=0; B1=0; B0=0; P3=0; P2=1; P1=1; P0=1;
	#1 V2=0; V1=0; V0=0; B2=0; B1=0; B0=0; P3=1; P2=0; P1=0; P0=0;	
	end 
	
  initial
    #50 $finish;
  initial begin
      $dumpfile("FSM_tb.vcd");
      $dumpvars(0, testbench);
    end
  endmodule
	
	
	
	
	
	
	
	
	